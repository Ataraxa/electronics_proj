library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fpga_toplvl_testbench is 
end entity fpga_toplvl_testbench;