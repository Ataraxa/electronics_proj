library IEEE;
use IEEE.std_logic_1164.all;

entity REPROG_LUT is 
    port (
        input : in std_logic_vector(3 downto 0);
        output : 
    )